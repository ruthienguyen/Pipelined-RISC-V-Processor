`timescale 1ns / 1ps

module and1
    (input logic  a,
     input logic b,
     output logic  y);


assign y = a & b;

endmodule
