`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2018 10:22:44 PM
// Design Name: 
// Module Name: imm_Gen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//    localparam R_TYPE = 7'b0110011;
//    localparam LW     = 7'b0000011; // done
//    localparam SW     = 7'b0100011; // done
//    localparam BR     = 7'b1100011; // done
//    localparam RTypeI = 7'b0010011; //addi,ori,andi // done
//    U_TYPE // done
//    J_TYPE // done
// Utype?

module imm_Gen(
    input logic [31:0] inst_code,
    output logic [31:0] Imm_out);


always_comb
    case(inst_code[6:0])
        
        /*Base types*/
        7'b0000011 /*I-type load*/     : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[31:20]};
        7'b1100111 /*I-type jalr*/     : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[31:20]};
        7'b0100011 /*S-type*/    : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[31:25], inst_code[11:7]};
        7'b1100011 /*B-type*/   :
            Imm_out = {inst_code[31]? 19'b1:19'b0 , inst_code[31], inst_code[7], inst_code[30:25], inst_code[11:8], 1'b0};
        7'b1101111 /*J-type*/   :
             Imm_out = {inst_code[31]? 11'b1:11'b0 , inst_code[31], inst_code[19:12], inst_code[20], inst_code[30:25], inst_code[24:21], 1'b0};
       
       /*U-type*/

        7'b0010111 /*U-type auipc*/   :
            Imm_out = {inst_code[31], inst_code[30:20], inst_code[19:12], 12'b0};
        7'b0110111 /*U-type I lui*/    : 
            Imm_out = {inst_code[31], inst_code[30:20], inst_code[19:12], 12'b0};
       
       /*Immediates*/
        7'b0010011 /*I-type I*/     : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[31:20]};  
       7'b0100011 /*J-type I*/    : 
            Imm_out = {inst_code[31]? 10'b1:10'b0 , inst_code[19:12], inst_code[20], inst_code[30:25], inst_code[24:21], 1'b0};
        7'b0100011 /*B-type I*/    : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[7], inst_code[30:25], inst[11:8],1'b0};
        7'b0100011 /*S-type I*/    : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[30:25], inst_code[11:8], inst[7]};
        7'b0010011 /*R-type I*/     : 
            Imm_out = {inst_code[31]? 20'b1:20'b0 , inst_code[31:20]};
        default                    : 
            Imm_out = {32'b0};
    endcase
    
endmodule
